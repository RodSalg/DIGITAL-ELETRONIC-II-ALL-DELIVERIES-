library verilog;
use verilog.vl_types.all;
entity schematic_vlg_vec_tst is
end schematic_vlg_vec_tst;
