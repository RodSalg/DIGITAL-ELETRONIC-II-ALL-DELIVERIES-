library verilog;
use verilog.vl_types.all;
entity lgc_h0_vlg_vec_tst is
end lgc_h0_vlg_vec_tst;
