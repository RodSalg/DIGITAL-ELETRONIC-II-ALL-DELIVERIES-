library verilog;
use verilog.vl_types.all;
entity dsf_timer_vlg_vec_tst is
end dsf_timer_vlg_vec_tst;
