library verilog;
use verilog.vl_types.all;
entity dsf_timer_vlg_check_tst is
    port(
        count           : in     vl_logic_vector(3 downto 0);
        q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end dsf_timer_vlg_check_tst;
