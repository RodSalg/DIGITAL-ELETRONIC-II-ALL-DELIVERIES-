library verilog;
use verilog.vl_types.all;
entity rlc_microservice_vlg_vec_tst is
end rlc_microservice_vlg_vec_tst;
