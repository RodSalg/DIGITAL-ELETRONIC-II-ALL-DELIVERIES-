-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Sat Feb 12 01:35:57 2022"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY dsff_freqdivider23 IS 
	PORT
	(
		enable :  IN  STD_LOGIC;
		reset :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		q :  OUT  STD_LOGIC;
		count :  OUT  STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END dsff_freqdivider23;

ARCHITECTURE bdf_type OF dsff_freqdivider23 IS 

COMPONENT dsf_freqdivider
	PORT(enable : IN STD_LOGIC;
		 areset : IN STD_LOGIC;
		 clk : IN STD_LOGIC;
		 q : OUT STD_LOGIC;
		 count : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END COMPONENT;



BEGIN 



b2v_inst : dsf_freqdivider
PORT MAP(enable => enable,
		 areset => reset,
		 clk => clk,
		 q => q,
		 count => count);


END bdf_type;