library verilog;
use verilog.vl_types.all;
entity radar_eletronico_vlg_vec_tst is
end radar_eletronico_vlg_vec_tst;
